// soc_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                           //                       clk.clk
		output wire        hps_hps_io_emac1_inst_TX_CLK,      //                       hps.hps_io_emac1_inst_TX_CLK
		output wire        hps_hps_io_emac1_inst_TXD0,        //                          .hps_io_emac1_inst_TXD0
		output wire        hps_hps_io_emac1_inst_TXD1,        //                          .hps_io_emac1_inst_TXD1
		output wire        hps_hps_io_emac1_inst_TXD2,        //                          .hps_io_emac1_inst_TXD2
		output wire        hps_hps_io_emac1_inst_TXD3,        //                          .hps_io_emac1_inst_TXD3
		input  wire        hps_hps_io_emac1_inst_RXD0,        //                          .hps_io_emac1_inst_RXD0
		inout  wire        hps_hps_io_emac1_inst_MDIO,        //                          .hps_io_emac1_inst_MDIO
		output wire        hps_hps_io_emac1_inst_MDC,         //                          .hps_io_emac1_inst_MDC
		input  wire        hps_hps_io_emac1_inst_RX_CTL,      //                          .hps_io_emac1_inst_RX_CTL
		output wire        hps_hps_io_emac1_inst_TX_CTL,      //                          .hps_io_emac1_inst_TX_CTL
		input  wire        hps_hps_io_emac1_inst_RX_CLK,      //                          .hps_io_emac1_inst_RX_CLK
		input  wire        hps_hps_io_emac1_inst_RXD1,        //                          .hps_io_emac1_inst_RXD1
		input  wire        hps_hps_io_emac1_inst_RXD2,        //                          .hps_io_emac1_inst_RXD2
		input  wire        hps_hps_io_emac1_inst_RXD3,        //                          .hps_io_emac1_inst_RXD3
		inout  wire        hps_hps_io_sdio_inst_CMD,          //                          .hps_io_sdio_inst_CMD
		inout  wire        hps_hps_io_sdio_inst_D0,           //                          .hps_io_sdio_inst_D0
		inout  wire        hps_hps_io_sdio_inst_D1,           //                          .hps_io_sdio_inst_D1
		output wire        hps_hps_io_sdio_inst_CLK,          //                          .hps_io_sdio_inst_CLK
		inout  wire        hps_hps_io_sdio_inst_D2,           //                          .hps_io_sdio_inst_D2
		inout  wire        hps_hps_io_sdio_inst_D3,           //                          .hps_io_sdio_inst_D3
		inout  wire        hps_hps_io_usb1_inst_D0,           //                          .hps_io_usb1_inst_D0
		inout  wire        hps_hps_io_usb1_inst_D1,           //                          .hps_io_usb1_inst_D1
		inout  wire        hps_hps_io_usb1_inst_D2,           //                          .hps_io_usb1_inst_D2
		inout  wire        hps_hps_io_usb1_inst_D3,           //                          .hps_io_usb1_inst_D3
		inout  wire        hps_hps_io_usb1_inst_D4,           //                          .hps_io_usb1_inst_D4
		inout  wire        hps_hps_io_usb1_inst_D5,           //                          .hps_io_usb1_inst_D5
		inout  wire        hps_hps_io_usb1_inst_D6,           //                          .hps_io_usb1_inst_D6
		inout  wire        hps_hps_io_usb1_inst_D7,           //                          .hps_io_usb1_inst_D7
		input  wire        hps_hps_io_usb1_inst_CLK,          //                          .hps_io_usb1_inst_CLK
		output wire        hps_hps_io_usb1_inst_STP,          //                          .hps_io_usb1_inst_STP
		input  wire        hps_hps_io_usb1_inst_DIR,          //                          .hps_io_usb1_inst_DIR
		input  wire        hps_hps_io_usb1_inst_NXT,          //                          .hps_io_usb1_inst_NXT
		output wire        hps_hps_io_spim1_inst_CLK,         //                          .hps_io_spim1_inst_CLK
		output wire        hps_hps_io_spim1_inst_MOSI,        //                          .hps_io_spim1_inst_MOSI
		input  wire        hps_hps_io_spim1_inst_MISO,        //                          .hps_io_spim1_inst_MISO
		output wire        hps_hps_io_spim1_inst_SS0,         //                          .hps_io_spim1_inst_SS0
		input  wire        hps_hps_io_uart0_inst_RX,          //                          .hps_io_uart0_inst_RX
		output wire        hps_hps_io_uart0_inst_TX,          //                          .hps_io_uart0_inst_TX
		inout  wire        hps_hps_io_i2c0_inst_SDA,          //                          .hps_io_i2c0_inst_SDA
		inout  wire        hps_hps_io_i2c0_inst_SCL,          //                          .hps_io_i2c0_inst_SCL
		inout  wire        hps_hps_io_i2c1_inst_SDA,          //                          .hps_io_i2c1_inst_SDA
		inout  wire        hps_hps_io_i2c1_inst_SCL,          //                          .hps_io_i2c1_inst_SCL
		inout  wire        hps_hps_io_gpio_inst_GPIO09,       //                          .hps_io_gpio_inst_GPIO09
		inout  wire        hps_hps_io_gpio_inst_GPIO35,       //                          .hps_io_gpio_inst_GPIO35
		inout  wire        hps_hps_io_gpio_inst_GPIO40,       //                          .hps_io_gpio_inst_GPIO40
		inout  wire        hps_hps_io_gpio_inst_GPIO48,       //                          .hps_io_gpio_inst_GPIO48
		inout  wire        hps_hps_io_gpio_inst_GPIO53,       //                          .hps_io_gpio_inst_GPIO53
		inout  wire        hps_hps_io_gpio_inst_GPIO54,       //                          .hps_io_gpio_inst_GPIO54
		inout  wire        hps_hps_io_gpio_inst_GPIO61,       //                          .hps_io_gpio_inst_GPIO61
		input  wire        hps_0_f2h_cold_reset_req_reset_n,  //  hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n, // hps_0_f2h_debug_reset_req.reset_n
		input  wire        hps_0_f2h_dma_req0_dma_req,        //        hps_0_f2h_dma_req0.dma_req
		input  wire        hps_0_f2h_dma_req0_dma_single,     //                          .dma_single
		output wire        hps_0_f2h_dma_req0_dma_ack,        //                          .dma_ack
		input  wire        hps_0_f2h_dma_req1_dma_req,        //        hps_0_f2h_dma_req1.dma_req
		input  wire        hps_0_f2h_dma_req1_dma_single,     //                          .dma_single
		output wire        hps_0_f2h_dma_req1_dma_ack,        //                          .dma_ack
		input  wire        hps_0_f2h_warm_reset_req_reset_n,  //  hps_0_f2h_warm_reset_req.reset_n
		output wire        hps_0_h2f_reset_reset_n,           //           hps_0_h2f_reset.reset_n
		output wire [14:0] hps_ddr3_mem_a,                    //                  hps_ddr3.mem_a
		output wire [2:0]  hps_ddr3_mem_ba,                   //                          .mem_ba
		output wire        hps_ddr3_mem_ck,                   //                          .mem_ck
		output wire        hps_ddr3_mem_ck_n,                 //                          .mem_ck_n
		output wire        hps_ddr3_mem_cke,                  //                          .mem_cke
		output wire        hps_ddr3_mem_cs_n,                 //                          .mem_cs_n
		output wire        hps_ddr3_mem_ras_n,                //                          .mem_ras_n
		output wire        hps_ddr3_mem_cas_n,                //                          .mem_cas_n
		output wire        hps_ddr3_mem_we_n,                 //                          .mem_we_n
		output wire        hps_ddr3_mem_reset_n,              //                          .mem_reset_n
		inout  wire [31:0] hps_ddr3_mem_dq,                   //                          .mem_dq
		inout  wire [3:0]  hps_ddr3_mem_dqs,                  //                          .mem_dqs
		inout  wire [3:0]  hps_ddr3_mem_dqs_n,                //                          .mem_dqs_n
		output wire        hps_ddr3_mem_odt,                  //                          .mem_odt
		output wire [3:0]  hps_ddr3_mem_dm,                   //                          .mem_dm
		input  wire        hps_ddr3_oct_rzqin,                //                          .oct_rzqin
		input  wire        loopback_fifo_0_rx_pri_ack,        //    loopback_fifo_0_rx_pri.ack
		output wire        loopback_fifo_0_rx_pri_burst,      //                          .burst
		output wire        loopback_fifo_0_rx_pri_single,     //                          .single
		output wire        loopback_fifo_0_tx_pri_single,     //    loopback_fifo_0_tx_pri.single
		input  wire        loopback_fifo_0_tx_pri_ack,        //                          .ack
		output wire        loopback_fifo_0_tx_pri_burst,      //                          .burst
		input  wire        reset_reset_n                      //                     reset.reset_n
	);

	wire   [1:0] hps_0_h2f_axi_master_awburst;                      // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                        // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [7:0] hps_0_h2f_axi_master_wstrb;                        // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                       // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                          // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                       // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                        // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                          // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                      // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                       // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                       // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                       // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                       // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [63:0] hps_0_h2f_axi_master_wdata;                        // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                      // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                      // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                         // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                       // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                       // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                       // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                        // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                      // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [63:0] hps_0_h2f_axi_master_rdata;                        // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                      // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                      // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                       // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                       // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                        // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                        // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                        // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                         // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                          // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                       // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                       // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                      // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                       // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire  [63:0] mm_interconnect_0_loopback_fifo_0_data_readdata;   // Loopback_FIFO_0:d_readdata -> mm_interconnect_0:Loopback_FIFO_0_data_readdata
	wire   [0:0] mm_interconnect_0_loopback_fifo_0_data_address;    // mm_interconnect_0:Loopback_FIFO_0_data_address -> Loopback_FIFO_0:d_address
	wire         mm_interconnect_0_loopback_fifo_0_data_read;       // mm_interconnect_0:Loopback_FIFO_0_data_read -> Loopback_FIFO_0:d_read
	wire   [7:0] mm_interconnect_0_loopback_fifo_0_data_byteenable; // mm_interconnect_0:Loopback_FIFO_0_data_byteenable -> Loopback_FIFO_0:d_byteenable
	wire         mm_interconnect_0_loopback_fifo_0_data_write;      // mm_interconnect_0:Loopback_FIFO_0_data_write -> Loopback_FIFO_0:d_write
	wire  [63:0] mm_interconnect_0_loopback_fifo_0_data_writedata;  // mm_interconnect_0:Loopback_FIFO_0_data_writedata -> Loopback_FIFO_0:d_writedata
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                   // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                     // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                     // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                    // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                    // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                     // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                       // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                   // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                    // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                    // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                    // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                    // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                     // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                   // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                   // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                      // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                    // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                    // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                    // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                     // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                   // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                     // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                   // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                   // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                    // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                    // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                     // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                     // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                     // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                      // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                    // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                    // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                   // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                    // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_1_loopback_fifo_0_csr_readdata;    // Loopback_FIFO_0:csr_readdata -> mm_interconnect_1:Loopback_FIFO_0_csr_readdata
	wire   [2:0] mm_interconnect_1_loopback_fifo_0_csr_address;     // mm_interconnect_1:Loopback_FIFO_0_csr_address -> Loopback_FIFO_0:csr_address
	wire         mm_interconnect_1_loopback_fifo_0_csr_read;        // mm_interconnect_1:Loopback_FIFO_0_csr_read -> Loopback_FIFO_0:csr_read
	wire   [3:0] mm_interconnect_1_loopback_fifo_0_csr_byteenable;  // mm_interconnect_1:Loopback_FIFO_0_csr_byteenable -> Loopback_FIFO_0:csr_byteenable
	wire         mm_interconnect_1_loopback_fifo_0_csr_write;       // mm_interconnect_1:Loopback_FIFO_0_csr_write -> Loopback_FIFO_0:csr_write
	wire  [31:0] mm_interconnect_1_loopback_fifo_0_csr_writedata;   // mm_interconnect_1:Loopback_FIFO_0_csr_writedata -> Loopback_FIFO_0:csr_writedata
	wire  [31:0] hps_0_f2h_irq0_irq;                                // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                    // rst_controller:reset_out -> [Loopback_FIFO_0:reset, mm_interconnect_0:Loopback_FIFO_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:Loopback_FIFO_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                // rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	flow_control_fifo #(
		.DATA_WIDTH (64),
		.FIFO_DEPTH (1024)
	) loopback_fifo_0 (
		.clk            (clk_clk),                                           //  clock.clk
		.reset          (rst_controller_reset_out_reset),                    //  reset.reset
		.csr_address    (mm_interconnect_1_loopback_fifo_0_csr_address),     //    csr.address
		.csr_write      (mm_interconnect_1_loopback_fifo_0_csr_write),       //       .write
		.csr_writedata  (mm_interconnect_1_loopback_fifo_0_csr_writedata),   //       .writedata
		.csr_byteenable (mm_interconnect_1_loopback_fifo_0_csr_byteenable),  //       .byteenable
		.csr_read       (mm_interconnect_1_loopback_fifo_0_csr_read),        //       .read
		.csr_readdata   (mm_interconnect_1_loopback_fifo_0_csr_readdata),    //       .readdata
		.d_address      (mm_interconnect_0_loopback_fifo_0_data_address),    //   data.address
		.d_write        (mm_interconnect_0_loopback_fifo_0_data_write),      //       .write
		.d_writedata    (mm_interconnect_0_loopback_fifo_0_data_writedata),  //       .writedata
		.d_byteenable   (mm_interconnect_0_loopback_fifo_0_data_byteenable), //       .byteenable
		.d_read         (mm_interconnect_0_loopback_fifo_0_data_read),       //       .read
		.d_readdata     (mm_interconnect_0_loopback_fifo_0_data_readdata),   //       .readdata
		.tx_single      (loopback_fifo_0_tx_pri_single),                     // tx_pri.single
		.tx_ack         (loopback_fifo_0_tx_pri_ack),                        //       .ack
		.tx_burst       (loopback_fifo_0_tx_pri_burst),                      //       .burst
		.rx_ack         (loopback_fifo_0_rx_pri_ack),                        // rx_pri.ack
		.rx_burst       (loopback_fifo_0_rx_pri_burst),                      //       .burst
		.rx_single      (loopback_fifo_0_rx_pri_single)                      //       .single
	);

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),  //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n), // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),  //  f2h_warm_reset_req.reset_n
		.h2f_user1_clk            (),                                  //     h2f_user1_clock.clk
		.f2h_dma_req0_req         (hps_0_f2h_dma_req0_dma_req),        //        f2h_dma_req0.dma_req
		.f2h_dma_req0_single      (hps_0_f2h_dma_req0_dma_single),     //                    .dma_single
		.f2h_dma_req0_ack         (hps_0_f2h_dma_req0_dma_ack),        //                    .dma_ack
		.f2h_dma_req1_req         (hps_0_f2h_dma_req1_dma_req),        //        f2h_dma_req1.dma_req
		.f2h_dma_req1_single      (hps_0_f2h_dma_req1_dma_single),     //                    .dma_single
		.f2h_dma_req1_ack         (hps_0_f2h_dma_req1_dma_ack),        //                    .dma_ack
		.mem_a                    (hps_ddr3_mem_a),                    //              memory.mem_a
		.mem_ba                   (hps_ddr3_mem_ba),                   //                    .mem_ba
		.mem_ck                   (hps_ddr3_mem_ck),                   //                    .mem_ck
		.mem_ck_n                 (hps_ddr3_mem_ck_n),                 //                    .mem_ck_n
		.mem_cke                  (hps_ddr3_mem_cke),                  //                    .mem_cke
		.mem_cs_n                 (hps_ddr3_mem_cs_n),                 //                    .mem_cs_n
		.mem_ras_n                (hps_ddr3_mem_ras_n),                //                    .mem_ras_n
		.mem_cas_n                (hps_ddr3_mem_cas_n),                //                    .mem_cas_n
		.mem_we_n                 (hps_ddr3_mem_we_n),                 //                    .mem_we_n
		.mem_reset_n              (hps_ddr3_mem_reset_n),              //                    .mem_reset_n
		.mem_dq                   (hps_ddr3_mem_dq),                   //                    .mem_dq
		.mem_dqs                  (hps_ddr3_mem_dqs),                  //                    .mem_dqs
		.mem_dqs_n                (hps_ddr3_mem_dqs_n),                //                    .mem_dqs_n
		.mem_odt                  (hps_ddr3_mem_odt),                  //                    .mem_odt
		.mem_dm                   (hps_ddr3_mem_dm),                   //                    .mem_dm
		.oct_rzqin                (hps_ddr3_oct_rzqin),                //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_hps_io_emac1_inst_TX_CLK),      //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_hps_io_emac1_inst_TXD0),        //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_hps_io_emac1_inst_TXD1),        //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_hps_io_emac1_inst_TXD2),        //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_hps_io_emac1_inst_TXD3),        //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_hps_io_emac1_inst_RXD0),        //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_hps_io_emac1_inst_MDIO),        //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_hps_io_emac1_inst_MDC),         //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_hps_io_emac1_inst_RX_CTL),      //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_hps_io_emac1_inst_TX_CTL),      //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_hps_io_emac1_inst_RX_CLK),      //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_hps_io_emac1_inst_RXD1),        //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_hps_io_emac1_inst_RXD2),        //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_hps_io_emac1_inst_RXD3),        //                    .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_hps_io_sdio_inst_CMD),          //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_hps_io_sdio_inst_D0),           //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_hps_io_sdio_inst_D1),           //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_hps_io_sdio_inst_CLK),          //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_hps_io_sdio_inst_D2),           //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_hps_io_sdio_inst_D3),           //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_hps_io_usb1_inst_D0),           //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_hps_io_usb1_inst_D1),           //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_hps_io_usb1_inst_D2),           //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_hps_io_usb1_inst_D3),           //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_hps_io_usb1_inst_D4),           //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_hps_io_usb1_inst_D5),           //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_hps_io_usb1_inst_D6),           //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_hps_io_usb1_inst_D7),           //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_hps_io_usb1_inst_CLK),          //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_hps_io_usb1_inst_STP),          //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_hps_io_usb1_inst_DIR),          //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_hps_io_usb1_inst_NXT),          //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_hps_io_spim1_inst_CLK),         //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_hps_io_spim1_inst_MOSI),        //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_hps_io_spim1_inst_MISO),        //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_hps_io_spim1_inst_SS0),         //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_hps_io_uart0_inst_RX),          //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_hps_io_uart0_inst_TX),          //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_hps_io_i2c0_inst_SDA),          //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_hps_io_i2c0_inst_SCL),          //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_hps_io_i2c1_inst_SDA),          //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_hps_io_i2c1_inst_SCL),          //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_hps_io_gpio_inst_GPIO09),       //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_hps_io_gpio_inst_GPIO35),       //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_hps_io_gpio_inst_GPIO40),       //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_hps_io_gpio_inst_GPIO48),       //                    .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_hps_io_gpio_inst_GPIO53),       //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_hps_io_gpio_inst_GPIO54),       //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_hps_io_gpio_inst_GPIO61),       //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),           //           h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                           //       h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),         //      h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),       //                    .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),        //                    .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),       //                    .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),      //                    .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),       //                    .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),      //                    .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),       //                    .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),      //                    .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),      //                    .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),          //                    .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),        //                    .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),        //                    .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),        //                    .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),       //                    .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),       //                    .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),          //                    .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),        //                    .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),       //                    .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),       //                    .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),         //                    .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),       //                    .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),        //                    .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),       //                    .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),      //                    .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),       //                    .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),      //                    .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),       //                    .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),      //                    .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),      //                    .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),          //                    .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),        //                    .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),        //                    .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),        //                    .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),       //                    .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),       //                    .rready
		.f2h_axi_clk              (clk_clk),                           //       f2h_axi_clock.clk
		.f2h_AWID                 (),                                  //       f2h_axi_slave.awid
		.f2h_AWADDR               (),                                  //                    .awaddr
		.f2h_AWLEN                (),                                  //                    .awlen
		.f2h_AWSIZE               (),                                  //                    .awsize
		.f2h_AWBURST              (),                                  //                    .awburst
		.f2h_AWLOCK               (),                                  //                    .awlock
		.f2h_AWCACHE              (),                                  //                    .awcache
		.f2h_AWPROT               (),                                  //                    .awprot
		.f2h_AWVALID              (),                                  //                    .awvalid
		.f2h_AWREADY              (),                                  //                    .awready
		.f2h_AWUSER               (),                                  //                    .awuser
		.f2h_WID                  (),                                  //                    .wid
		.f2h_WDATA                (),                                  //                    .wdata
		.f2h_WSTRB                (),                                  //                    .wstrb
		.f2h_WLAST                (),                                  //                    .wlast
		.f2h_WVALID               (),                                  //                    .wvalid
		.f2h_WREADY               (),                                  //                    .wready
		.f2h_BID                  (),                                  //                    .bid
		.f2h_BRESP                (),                                  //                    .bresp
		.f2h_BVALID               (),                                  //                    .bvalid
		.f2h_BREADY               (),                                  //                    .bready
		.f2h_ARID                 (),                                  //                    .arid
		.f2h_ARADDR               (),                                  //                    .araddr
		.f2h_ARLEN                (),                                  //                    .arlen
		.f2h_ARSIZE               (),                                  //                    .arsize
		.f2h_ARBURST              (),                                  //                    .arburst
		.f2h_ARLOCK               (),                                  //                    .arlock
		.f2h_ARCACHE              (),                                  //                    .arcache
		.f2h_ARPROT               (),                                  //                    .arprot
		.f2h_ARVALID              (),                                  //                    .arvalid
		.f2h_ARREADY              (),                                  //                    .arready
		.f2h_ARUSER               (),                                  //                    .aruser
		.f2h_RID                  (),                                  //                    .rid
		.f2h_RDATA                (),                                  //                    .rdata
		.f2h_RRESP                (),                                  //                    .rresp
		.f2h_RLAST                (),                                  //                    .rlast
		.f2h_RVALID               (),                                  //                    .rvalid
		.f2h_RREADY               (),                                  //                    .rready
		.h2f_lw_axi_clk           (clk_clk),                           //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),      //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),    //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),     //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),    //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),   //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),    //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),   //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),    //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),   //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),   //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),       //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),     //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),     //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),     //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),    //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),    //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),       //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),     //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),    //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),    //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),      //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),    //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),     //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),    //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),   //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),    //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),   //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),    //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),   //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),   //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),       //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),     //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),     //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),     //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),    //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),    //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                 //            f2h_irq1.irq
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                         //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                       //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                        //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                       //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                      //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                       //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                      //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                       //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                      //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                      //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                          //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                        //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                        //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                        //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                       //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                       //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                          //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                        //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                       //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                       //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                         //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                       //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                        //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                       //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                      //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                       //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                      //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                       //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                      //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                      //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                          //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                        //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                        //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                        //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                       //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                       //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                           //                                                  clk_0_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.Loopback_FIFO_0_reset_reset_bridge_in_reset_reset                (rst_controller_reset_out_reset),                    //                Loopback_FIFO_0_reset_reset_bridge_in_reset.reset
		.Loopback_FIFO_0_data_address                                     (mm_interconnect_0_loopback_fifo_0_data_address),    //                                       Loopback_FIFO_0_data.address
		.Loopback_FIFO_0_data_write                                       (mm_interconnect_0_loopback_fifo_0_data_write),      //                                                           .write
		.Loopback_FIFO_0_data_read                                        (mm_interconnect_0_loopback_fifo_0_data_read),       //                                                           .read
		.Loopback_FIFO_0_data_readdata                                    (mm_interconnect_0_loopback_fifo_0_data_readdata),   //                                                           .readdata
		.Loopback_FIFO_0_data_writedata                                   (mm_interconnect_0_loopback_fifo_0_data_writedata),  //                                                           .writedata
		.Loopback_FIFO_0_data_byteenable                                  (mm_interconnect_0_loopback_fifo_0_data_byteenable)  //                                                           .byteenable
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                     //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                   //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                    //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                   //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                  //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                   //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                  //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                   //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                  //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                  //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                      //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                    //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                    //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                    //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                   //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                   //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                      //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                    //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                   //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                   //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                     //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                   //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                    //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                   //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                  //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                   //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                  //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                   //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                  //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                  //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                      //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                    //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                    //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                    //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                   //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                   //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                          //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),               // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.Loopback_FIFO_0_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                   //                   Loopback_FIFO_0_reset_reset_bridge_in_reset.reset
		.Loopback_FIFO_0_csr_address                                         (mm_interconnect_1_loopback_fifo_0_csr_address),    //                                           Loopback_FIFO_0_csr.address
		.Loopback_FIFO_0_csr_write                                           (mm_interconnect_1_loopback_fifo_0_csr_write),      //                                                              .write
		.Loopback_FIFO_0_csr_read                                            (mm_interconnect_1_loopback_fifo_0_csr_read),       //                                                              .read
		.Loopback_FIFO_0_csr_readdata                                        (mm_interconnect_1_loopback_fifo_0_csr_readdata),   //                                                              .readdata
		.Loopback_FIFO_0_csr_writedata                                       (mm_interconnect_1_loopback_fifo_0_csr_writedata),  //                                                              .writedata
		.Loopback_FIFO_0_csr_byteenable                                      (mm_interconnect_1_loopback_fifo_0_csr_byteenable)  //                                                              .byteenable
	);

	soc_system_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
